library verilog;
use verilog.vl_types.all;
entity Tx_TB is
end Tx_TB;
