library verilog;
use verilog.vl_types.all;
entity ripple_counter_TB is
end ripple_counter_TB;
