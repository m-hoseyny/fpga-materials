library verilog;
use verilog.vl_types.all;
entity tb_Rx is
end tb_Rx;
