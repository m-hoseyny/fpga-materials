library verilog;
use verilog.vl_types.all;
entity test_overlap_nonoverlap is
end test_overlap_nonoverlap;
