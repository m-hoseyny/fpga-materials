library verilog;
use verilog.vl_types.all;
entity rx_tx_test is
end rx_tx_test;
