library verilog;
use verilog.vl_types.all;
entity Ram_TB is
end Ram_TB;
