library verilog;
use verilog.vl_types.all;
entity Mult_TB is
end Mult_TB;
