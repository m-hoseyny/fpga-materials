library verilog;
use verilog.vl_types.all;
entity CoeffRam_TB is
end CoeffRam_TB;
