library verilog;
use verilog.vl_types.all;
entity SE_TB is
end SE_TB;
