library verilog;
use verilog.vl_types.all;
entity BRG_TB is
end BRG_TB;
