library verilog;
use verilog.vl_types.all;
entity DI_TB is
end DI_TB;
