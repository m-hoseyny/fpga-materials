library verilog;
use verilog.vl_types.all;
entity Registe_TB is
end Registe_TB;
