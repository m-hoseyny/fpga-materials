library verilog;
use verilog.vl_types.all;
entity test_dut is
end test_dut;
