library verilog;
use verilog.vl_types.all;
entity Counter_TB is
end Counter_TB;
